module Teste(input  K, 
				output L);

	assign L= K;
	
endmodule
