module Display(input [3:0]E,
					output reg[0:6] S);
					
		always@(*)begin
	case(E)
		4'b0000:S=7'b0000001;
		4'b0001:S=7'b1001111;
		4'b0010:S=7'b0010010;
		4'b0011:S=7'b0000110;
		4'b0100:S=7'b1001100;
		4'b0101:S=7'b0100100;
		4'b0110:S=7'b0100000;
		4'b0111:S=7'b0001111;
		4'b1000:S=7'b0000000;
		4'b1001:S=7'b0001100;
		4'b1010:S=7'b0001000;
		4'b1011:S=7'b1100000;
		4'b1100:S=7'b0110001;
		4'b1101:S=7'b1000010;
		4'b1110:S=7'b0110000;
		4'b1111:S=7'b0111000;
	endcase
	end
endmodule
